
module ariane_Soc_Wrap (
	input sys_clk,
	input RSTn,
	
	input irq,


(* X_INTERFACE_PARAMETER = "FREQ_HZ 30000000" *)
    output wire [3 : 0] PERIP_AXI_AWID,
    output wire [63 : 0] PERIP_AXI_AWADDR,
    output wire [7 : 0] PERIP_AXI_AWLEN,
    output wire [2 : 0] PERIP_AXI_AWSIZE,
    output wire [1 : 0] PERIP_AXI_AWBURST,
    output wire PERIP_AXI_AWLOCK,
    output wire [3 : 0] PERIP_AXI_AWCACHE,
    output wire [2 : 0] PERIP_AXI_AWPROT,
    output wire PERIP_AXI_AWVALID,
    input wire  PERIP_AXI_AWREADY,
    output wire [63 : 0] PERIP_AXI_WDATA,
    output wire [7 : 0] PERIP_AXI_WSTRB,
    output wire PERIP_AXI_WLAST,
    output wire PERIP_AXI_WVALID,
    input wire PERIP_AXI_WREADY,
    input wire [3 : 0] PERIP_AXI_BID,
    input wire [1 : 0] PERIP_AXI_BRESP,
    input wire PERIP_AXI_BVALID,
    output wire PERIP_AXI_BREADY,
    output wire [3 : 0] PERIP_AXI_ARID,
    output wire [63 : 0] PERIP_AXI_ARADDR,
    output wire [7 : 0] PERIP_AXI_ARLEN,
    output wire [2 : 0] PERIP_AXI_ARSIZE,
    output wire [1 : 0] PERIP_AXI_ARBURST,
    output wire  PERIP_AXI_ARLOCK,
    output wire [3 : 0] PERIP_AXI_ARCACHE,
    output wire [2 : 0] PERIP_AXI_ARPROT,
    output wire  PERIP_AXI_ARVALID,
    input wire  PERIP_AXI_ARREADY,
    input wire [3 : 0] PERIP_AXI_RID,
    input wire [63 : 0] PERIP_AXI_RDATA,
    input wire [1 : 0] PERIP_AXI_RRESP,
    input wire PERIP_AXI_RLAST,
    input wire PERIP_AXI_RVALID,
    output wire PERIP_AXI_RREADY,
    output wire [4 : 0] PERIP_AXI_AWUSER,
    output wire [3 : 0] PERIP_AXI_AWQOS,
    output wire [4 : 0] PERIP_AXI_WUSER,
    input wire [4 : 0] PERIP_AXI_BUSER,
    output wire [4 : 0] PERIP_AXI_ARUSER,
    output wire [3 : 0] PERIP_AXI_ARQOS,
    input wire [4 : 0] PERIP_AXI_RUSER,
    output wire [3:0] PERIP_AXI_AWREGION,
    output wire [3:0] PERIP_AXI_ARREGION,


(* X_INTERFACE_PARAMETER = "FREQ_HZ 30000000" *)
	output wire [3 : 0] MEM_AXI_AWID,
	output wire [63 : 0] MEM_AXI_AWADDR,
	output wire [7 : 0] MEM_AXI_AWLEN,
	output wire [2 : 0] MEM_AXI_AWSIZE,
	output wire [1 : 0] MEM_AXI_AWBURST,
	output wire  MEM_AXI_AWLOCK,
	output wire [3 : 0] MEM_AXI_AWCACHE,
	output wire [2 : 0] MEM_AXI_AWPROT,
	// output wire [3 : 0] MEM_AXI_AWQOS,
// output wire [C_M_AXI_AWUSER_WIDTH-1 : 0] MEM_AXI_AWUSER,
	output wire  MEM_AXI_AWVALID,
	input wire  MEM_AXI_AWREADY,
	output wire [63 : 0] MEM_AXI_WDATA,
	output wire [7 : 0] MEM_AXI_WSTRB,
	output wire  MEM_AXI_WLAST,
// output wire [C_M_AXI_WUSER_WIDTH-1 : 0] MEM_AXI_WUSER,
	output wire  MEM_AXI_WVALID,
	input wire  MEM_AXI_WREADY,
	input wire [3 : 0] MEM_AXI_BID,
	input wire [1 : 0] MEM_AXI_BRESP,
// input wire [C_M_AXI_BUSER_WIDTH-1 : 0] MEM_AXI_BUSER,
	input wire  MEM_AXI_BVALID,
	output wire  MEM_AXI_BREADY,
	output wire [3 : 0] MEM_AXI_ARID,
	output wire [63 : 0] MEM_AXI_ARADDR,
	output wire [7 : 0] MEM_AXI_ARLEN,
	output wire [2 : 0] MEM_AXI_ARSIZE,
	output wire [1 : 0] MEM_AXI_ARBURST,
	output wire  MEM_AXI_ARLOCK,
	output wire [3 : 0] MEM_AXI_ARCACHE,
	output wire [2 : 0] MEM_AXI_ARPROT,
// 	output wire [3 : 0] MEM_AXI_ARQOS,
// output wire [C_M_AXI_ARUSER_WIDTH-1 : 0] MEM_AXI_ARUSER,
	output wire  MEM_AXI_ARVALID,
	input wire  MEM_AXI_ARREADY,
	input wire [3 : 0] MEM_AXI_RID,
	input wire [63 : 0] MEM_AXI_RDATA,
	input wire [1 : 0] MEM_AXI_RRESP,
	input wire  MEM_AXI_RLAST,
// input wire [C_M_AXI_RUSER_WIDTH-1 : 0] MEM_AXI_RUSER,
	input wire  MEM_AXI_RVALID,
	output wire  MEM_AXI_RREADY,



	// common part
	// input trst_n,
	input tck,
	input tms,
	input tdi,
	output tdo
	
);




ariane_xilinx bd_xilinx(
	.sys_clk(sys_clk),
	.RSTn(RSTn),

	.irq({irq,1'b0}),
	// .sw(sw),

    .PERIP_AXI_AWID(PERIP_AXI_AWID),
    .PERIP_AXI_AWADDR(PERIP_AXI_AWADDR),
    .PERIP_AXI_AWLEN(PERIP_AXI_AWLEN),
    .PERIP_AXI_AWSIZE(PERIP_AXI_AWSIZE),
    .PERIP_AXI_AWBURST(PERIP_AXI_AWBURST),
    .PERIP_AXI_AWLOCK(PERIP_AXI_AWLOCK),
    .PERIP_AXI_AWCACHE(PERIP_AXI_AWCACHE),
    .PERIP_AXI_AWPROT(PERIP_AXI_AWPROT),
    .PERIP_AXI_AWVALID(PERIP_AXI_AWVALID),
    .PERIP_AXI_AWREADY(PERIP_AXI_AWREADY),
    .PERIP_AXI_WDATA(PERIP_AXI_WDATA),
    .PERIP_AXI_WSTRB(PERIP_AXI_WSTRB),
    .PERIP_AXI_WLAST(PERIP_AXI_WLAST),
    .PERIP_AXI_WVALID(PERIP_AXI_WVALID),
    .PERIP_AXI_WREADY(PERIP_AXI_WREADY),
    .PERIP_AXI_BID(PERIP_AXI_BID),
    .PERIP_AXI_BRESP(PERIP_AXI_BRESP),
    .PERIP_AXI_BVALID(PERIP_AXI_BVALID),
    .PERIP_AXI_BREADY(PERIP_AXI_BREADY),
    .PERIP_AXI_ARID(PERIP_AXI_ARID),
    .PERIP_AXI_ARADDR(PERIP_AXI_ARADDR),
    .PERIP_AXI_ARLEN(PERIP_AXI_ARLEN),
    .PERIP_AXI_ARSIZE(PERIP_AXI_ARSIZE),
    .PERIP_AXI_ARBURST(PERIP_AXI_ARBURST),
    .PERIP_AXI_ARLOCK(PERIP_AXI_ARLOCK),
    .PERIP_AXI_ARCACHE(PERIP_AXI_ARCACHE),
    .PERIP_AXI_ARPROT(PERIP_AXI_ARPROT),
    .PERIP_AXI_ARVALID(PERIP_AXI_ARVALID),
    .PERIP_AXI_ARREADY(PERIP_AXI_ARREADY),
    .PERIP_AXI_RID(PERIP_AXI_RID),
    .PERIP_AXI_RDATA(PERIP_AXI_RDATA),
    .PERIP_AXI_RRESP(PERIP_AXI_RRESP),
    .PERIP_AXI_RLAST(PERIP_AXI_RLAST),
    .PERIP_AXI_RVALID(PERIP_AXI_RVALID),
    .PERIP_AXI_RREADY(PERIP_AXI_RREADY),
    .PERIP_AXI_AWUSER(PERIP_AXI_AWUSER),
    .PERIP_AXI_AWQOS(PERIP_AXI_AWQOS),
    .PERIP_AXI_WUSER(PERIP_AXI_WUSER),
    .PERIP_AXI_BUSER(PERIP_AXI_BUSER),
    .PERIP_AXI_ARUSER(PERIP_AXI_ARUSER),
    .PERIP_AXI_ARQOS(PERIP_AXI_ARQOS),
    .PERIP_AXI_RUSER(PERIP_AXI_RUSER),
    .PERIP_AXI_AWREGION(PERIP_AXI_AWREGION),
    .PERIP_AXI_ARREGION(PERIP_AXI_ARREGION),



	.MEM_AXI_AWID(MEM_AXI_AWID),
	.MEM_AXI_AWADDR(MEM_AXI_AWADDR),
	.MEM_AXI_AWLEN(MEM_AXI_AWLEN),
	.MEM_AXI_AWSIZE(MEM_AXI_AWSIZE),
	.MEM_AXI_AWBURST(MEM_AXI_AWBURST),
	.MEM_AXI_AWLOCK(MEM_AXI_AWLOCK),
	.MEM_AXI_AWCACHE(MEM_AXI_AWCACHE),
	.MEM_AXI_AWPROT(MEM_AXI_AWPROT),
	.MEM_AXI_AWVALID(MEM_AXI_AWVALID),
	.MEM_AXI_AWREADY(MEM_AXI_AWREADY),
	.MEM_AXI_WDATA(MEM_AXI_WDATA),
	.MEM_AXI_WSTRB(MEM_AXI_WSTRB),
	.MEM_AXI_WLAST(MEM_AXI_WLAST),

	.MEM_AXI_WVALID(MEM_AXI_WVALID),
	.MEM_AXI_WREADY(MEM_AXI_WREADY),
	.MEM_AXI_BID(MEM_AXI_BID),
	.MEM_AXI_BRESP(MEM_AXI_BRESP),

	.MEM_AXI_BVALID(MEM_AXI_BVALID),
	.MEM_AXI_BREADY(MEM_AXI_BREADY),
	.MEM_AXI_ARID(MEM_AXI_ARID),
	.MEM_AXI_ARADDR(MEM_AXI_ARADDR),
	.MEM_AXI_ARLEN(MEM_AXI_ARLEN),
	.MEM_AXI_ARSIZE(MEM_AXI_ARSIZE),
	.MEM_AXI_ARBURST(MEM_AXI_ARBURST),
	.MEM_AXI_ARLOCK(MEM_AXI_ARLOCK),
	.MEM_AXI_ARCACHE(MEM_AXI_ARCACHE),
	.MEM_AXI_ARPROT(MEM_AXI_ARPROT),

	.MEM_AXI_ARVALID(MEM_AXI_ARVALID),
	.MEM_AXI_ARREADY(MEM_AXI_ARREADY),
	.MEM_AXI_RID(MEM_AXI_RID),
	.MEM_AXI_RDATA(MEM_AXI_RDATA),
	.MEM_AXI_RRESP(MEM_AXI_RRESP),
	.MEM_AXI_RLAST(MEM_AXI_RLAST),
	.MEM_AXI_RVALID(MEM_AXI_RVALID),
	.MEM_AXI_RREADY(MEM_AXI_RREADY),

	// common part
	// input trst_n,
	.tck(tck),
	.tms(tms),
	.tdi(tdi),
	.tdo(tdo)
);












endmodule


